`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Dexter Elmendorf
// Class:
// ECE 483 Lab #4
//
// Create Date: 06/16/2022
// File Name: Write_Decode.v
//
// Decoder for Write load into the Register Bank
//////////////////////////////////////////////////////////////////////////////////


module Write_Decode(
    input [4:0]RegAddr,
    input regWrite,
    
    output reg [31:0] regLoad
    );
   //Case each write address and set each corresponding load high
    always @(RegAddr, regWrite)
        case(RegAddr)
            5'b00000:regLoad <= 32'b00000000_00000000_00000000_00000001;
            5'b00001:regLoad <= 32'b00000000_00000000_00000000_00000010;
            5'b00010:regLoad <= 32'b00000000_00000000_00000000_00000100;
            5'b00011:regLoad <= 32'b00000000_00000000_00000000_00001000;
            5'b00100:regLoad <= 32'b00000000_00000000_00000000_00010000;
            5'b00101:regLoad <= 32'b00000000_00000000_00000000_00100000;
            5'b00110:regLoad <= 32'b00000000_00000000_00000000_01000000;
            5'b00111:regLoad <= 32'b00000000_00000000_00000000_10000000;
            5'b01000:regLoad <= 32'b00000000_00000000_00000001_00000000;
            5'b01001:regLoad <= 32'b00000000_00000000_00000010_00000000;
            5'b01010:regLoad <= 32'b00000000_00000000_00000100_00000000;
            5'b01011:regLoad <= 32'b00000000_00000000_00001000_00000000;
            5'b01100:regLoad <= 32'b00000000_00000000_00010000_00000000;
            5'b01101:regLoad <= 32'b00000000_00000000_00100000_00000000;
            5'b01110:regLoad <= 32'b00000000_00000000_01000000_00000000;
            5'b01111:regLoad <= 32'b00000000_00000000_10000000_00000000;
            5'b10000:regLoad <= 32'b00000000_00000001_00000000_00000000;
            5'b10001:regLoad <= 32'b00000000_00000010_00000000_00000000;
            5'b10010:regLoad <= 32'b00000000_00000100_00000000_00000000;
            5'b10011:regLoad <= 32'b00000000_00001000_00000000_00000000;
            5'b10100:regLoad <= 32'b00000000_00010000_00000000_00000000;
            5'b10101:regLoad <= 32'b00000000_00100000_00000000_00000000;
            5'b10110:regLoad <= 32'b00000000_01000000_00000000_00000000;
            5'b10111:regLoad <= 32'b00000000_10000000_00000000_00000000;
            5'b11000:regLoad <= 32'b00000001_00000000_00000000_00000000;
            5'b11001:regLoad <= 32'b00000010_00000000_00000000_00000000;
            5'b11010:regLoad <= 32'b00000100_00000000_00000000_00000000;
            5'b11011:regLoad <= 32'b00001000_00000000_00000000_00000000;
            5'b11100:regLoad <= 32'b00010000_00000000_00000000_00000000;
            5'b11101:regLoad <= 32'b00100000_00000000_00000000_00000000;
            5'b11110:regLoad <= 32'b01000000_00000000_00000000_00000000;
            5'b11111:regLoad <= 32'b10000000_00000000_00000000_00000000;
        endcase
endmodule