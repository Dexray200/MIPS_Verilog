`timescale 1ns / 1ps


module IR_Mem(output reg [31:0] data_out, input [31:0] address);
always@(address)begin
	case(address) 
	   // Program #1
	   /*
        32'h0000_0004: data_out = 32'b000000_00010_00011_00001_00000_100000;
        32'h0000_0008: data_out = 32'b000000_00101_00110_00100_00000_100010;
        32'h0000_000c: data_out = 32'b000000_01000_01001_00111_00000_100100;
        32'h0000_0010: data_out = 32'b000000_00001_01100_01010_00000_100101;
        32'h0000_0014: data_out = 32'b000000_00100_10001_10000_00000_101010;
        */
        
        //Program #2
        32'h0000_0004: data_out = 32'b000000_00011_00011_00001_00000_100000;
        32'h0000_0008: data_out = 32'b101011_00000_00010_00010_00000_010000;
        32'h0000_000c: data_out = 32'b000000_00001_00100_00111_00000_100100;
        32'h0000_0010: data_out = 32'b100011_00001_00111_00100_00000_000000;
        32'h0000_0014: data_out = 32'b100011_00101_00110_10000_00000_000110;   
        
        
		default: #7 data_out=32'h1234abcd;
	endcase
end

endmodule
